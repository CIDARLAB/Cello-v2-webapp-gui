module xor_gate(output out, input a, b);

   xor(out, a, b);

endmodule
