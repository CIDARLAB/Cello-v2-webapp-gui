module and_gate(output out, input a, b);

   and(out, a, b);

endmodule
